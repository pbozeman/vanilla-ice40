`ifndef DIRECTIVES_V
`define DIRECTIVES_V

// for simulation
`timescale 1ns / 1ps

// avoid undeclared symbols
`default_nettype none

`endif
