`timescale 1ns / 1ps


// pin 1 & 2 are the user LEDs.
// pin 21 is the clock. Skip those.

module solder_chk_top (
    input  wire clk_i,
    output wire led1_o,
    output wire led2_o,

    inout wire PIN3,
    inout wire PIN4,
    inout wire PIN7,
    inout wire PIN8,
    inout wire PIN9,
    inout wire PIN10,
    inout wire PIN11,
    inout wire PIN12,
    inout wire PIN15,
    inout wire PIN16,
    inout wire PIN17,
    inout wire PIN18,
    inout wire PIN19,
    inout wire PIN20,
    inout wire PIN22,
    inout wire PIN23,
    inout wire PIN24,
    inout wire PIN25,
    inout wire PIN26,
    inout wire PIN28,
    inout wire PIN29,
    inout wire PIN31,
    inout wire PIN32,
    inout wire PIN33,
    inout wire PIN34,
    inout wire PIN37,
    inout wire PIN38,
    inout wire PIN39,
    inout wire PIN41,
    inout wire PIN42,
    inout wire PIN43,
    inout wire PIN44,
    inout wire PIN45,
    inout wire PIN47,
    inout wire PIN48,
    inout wire PIN49,
    inout wire PIN52,
    inout wire PIN55,
    inout wire PIN56,
    inout wire PIN60,
    inout wire PIN61,
    inout wire PIN62,
    inout wire PIN63,
    inout wire PIN64,
    inout wire PIN67,
    inout wire PIN68,
    inout wire PIN70,
    inout wire PIN71,
    inout wire PIN73,
    inout wire PIN74,
    inout wire PIN75,
    inout wire PIN76,
    inout wire PIN78,
    inout wire PIN79,
    inout wire PIN80,
    inout wire PIN81,
    inout wire PIN82,
    inout wire PIN83,
    inout wire PIN84,
    inout wire PIN85,
    inout wire PIN87,
    inout wire PIN88,
    inout wire PIN90,
    inout wire PIN91,
    inout wire PIN93,
    inout wire PIN94,
    inout wire PIN95,
    inout wire PIN96,
    inout wire PIN97,
    inout wire PIN98,
    inout wire PIN99,
    inout wire PIN101,
    inout wire PIN102,
    inout wire PIN104,
    inout wire PIN105,
    inout wire PIN106,
    inout wire PIN107,
    inout wire PIN110,
    inout wire PIN112,
    inout wire PIN113,
    inout wire PIN114,
    inout wire PIN115,
    inout wire PIN116,
    inout wire PIN117,
    inout wire PIN118,
    inout wire PIN119,
    inout wire PIN120,
    inout wire PIN121,
    input wire PIN122,
    inout wire PIN124,
    inout wire PIN125,
    inout wire PIN128,
    inout wire PIN129,
    inout wire PIN130,
    inout wire PIN134,
    inout wire PIN135,
    inout wire PIN136,
    inout wire PIN137,
    inout wire PIN138,
    inout wire PIN139,
    inout wire PIN141,
    inout wire PIN142,
    inout wire PIN143,
    inout wire PIN144
);

  localparam NUM_PINS = 104;

  wire [NUM_PINS-1:0] test_pins;
  wire [NUM_PINS-1:0] result_pins;
  wire error;

  assign result_pins = {
    PIN3,
    PIN4,
    PIN7,
    PIN8,
    PIN9,
    PIN10,
    PIN11,
    PIN12,
    PIN15,
    PIN16,
    PIN17,
    PIN18,
    PIN19,
    PIN20,
    PIN22,
    PIN23,
    PIN24,
    PIN25,
    PIN26,
    PIN28,
    PIN29,
    PIN31,
    PIN32,
    PIN33,
    PIN34,
    PIN37,
    PIN38,
    PIN39,
    PIN41,
    PIN42,
    PIN43,
    PIN44,
    PIN45,
    PIN47,
    PIN48,
    PIN49,
    PIN52,
    PIN55,
    PIN56,
    PIN60,
    PIN61,
    PIN62,
    PIN63,
    PIN64,
    PIN67,
    PIN68,
    PIN70,
    PIN71,
    PIN73,
    PIN74,
    PIN75,
    PIN76,
    PIN78,
    PIN79,
    PIN80,
    PIN81,
    PIN82,
    PIN83,
    PIN84,
    PIN85,
    PIN87,
    PIN88,
    PIN90,
    PIN91,
    PIN93,
    PIN94,
    PIN95,
    PIN96,
    PIN97,
    PIN98,
    PIN99,
    PIN101,
    PIN102,
    PIN104,
    PIN105,
    PIN106,
    PIN107,
    PIN110,
    PIN112,
    PIN113,
    PIN114,
    PIN115,
    PIN116,
    PIN117,
    PIN118,
    PIN119,
    PIN120,
    PIN121,
    // PIN122,
    PIN124,
    PIN125,
    PIN128,
    PIN129,
    PIN130,
    PIN134,
    PIN135,
    PIN136,
    PIN137,
    PIN138,
    PIN139,
    PIN141,
    PIN142,
    PIN143,
    PIN144
  };

  assign {
    PIN3,
    PIN4,
    PIN7,
    PIN8,
    PIN9,
    PIN10,
    PIN11,
    PIN12,
    PIN15,
    PIN16,
    PIN17,
    PIN18,
    PIN19,
    PIN20,
    PIN22,
    PIN23,
    PIN24,
    PIN25,
    PIN26,
    PIN28,
    PIN29,
    PIN31,
    PIN32,
    PIN33,
    PIN34,
    PIN37,
    PIN38,
    PIN39,
    PIN41,
    PIN42,
    PIN43,
    PIN44,
    PIN45,
    PIN47,
    PIN48,
    PIN49,
    PIN52,
    PIN55,
    PIN56,
    PIN60,
    PIN61,
    PIN62,
    PIN63,
    PIN64,
    PIN67,
    PIN68,
    PIN70,
    PIN71,
    PIN73,
    PIN74,
    PIN75,
    PIN76,
    PIN78,
    PIN79,
    PIN80,
    PIN81,
    PIN82,
    PIN83,
    PIN84,
    PIN85,
    PIN87,
    PIN88,
    PIN90,
    PIN91,
    PIN93,
    PIN94,
    PIN95,
    PIN96,
    PIN97,
    PIN98,
    PIN99,
    PIN101,
    PIN102,
    PIN104,
    PIN105,
    PIN106,
    PIN107,
    PIN110,
    PIN112,
    PIN113,
    PIN114,
    PIN115,
    PIN116,
    PIN117,
    PIN118,
    PIN119,
    PIN120,
    PIN121,
    // PIN122,
    PIN124,
    PIN125,
    PIN128,
    PIN129,
    PIN130,
    PIN134,
    PIN135,
    PIN136,
    PIN137,
    PIN138,
    PIN139,
    PIN141,
    PIN142,
    PIN143,
    PIN144 } = test_pins;

  io_walker #(
      .NUM_PINS(103)
  ) uut (
      .clk_i(clk_i),
      .test_pins(test_pins),
      .result_pins(result_pins),
      .error_o(error)
  );

  assign led1_o = PIN122;
  assign led2_o = error;

endmodule
